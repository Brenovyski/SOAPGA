library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity soapga is
    port(
        clock        : in std_logic;
        reset        : in std_logic;
        ligar        : in std_logic;
        echo2        : in std_logic;
        echo1        : in std_logic;
        pwm          : out std_logic;
        trigger2     : out std_logic;
        trigger1     : out std_logic;
        saida_serial : out std_logic;
        sseg1        : out std_logic_vector(6 downto 0);
        sseg2        : out std_logic_vector(6 downto 0);
        sseg3        : out std_logic_vector(6 downto 0);
        sseg4        : out std_logic_vector(6 downto 0);
        db_estado    : out std_logic_vector(6 downto 0)
    );
end entity;

architecture soapga_arch of soapga is

    component soapga_uc is 
        port ( 
            clock            : in  std_logic;
            reset            : in  std_logic;
            ligar            : in  std_logic;
            pronto_medir1    : in  std_logic;
            pronto_medir2    : in  std_logic;
            mao_presente     : in  std_logic;
            fim_timer1       : in  std_logic;
            fim_timer2       : in  std_logic;
            pronto_tx        : in  std_logic;
            zera             : out std_logic;
            medir1           : out std_logic;
            medir2           : out std_logic;
            zera_timer1      : out std_logic;
            zera_timer2      : out std_logic;
            zera_hc          : out std_logic;
            conta_timer1     : out std_logic;
            conta_timer2     : out std_logic;
            gira_servo       : out std_logic;
            partida_tx       : out std_logic;
            sel              : out std_logic_vector(1 downto 0); 
            db_estado        : out std_logic_vector(3 downto 0)
        );
    end component;

    component soapga_fd is
        port (
            clock         : in std_logic;
            reset         : in std_logic;
            gira_servo    : in std_logic;
            medir2        : in std_logic;
            medir1        : in std_logic;
            echo2         : in std_logic;
            echo1         : in std_logic;
            sel           : in std_logic_vector(1 downto 0);
            partida_tx    : in std_logic;
            zera_timer1   : in std_logic;
            zera_timer2   : in std_logic;
            zera_hc       : in std_logic;
            conta_timer1  : in std_logic;
            conta_timer2  : in std_logic;
            pwm           : out std_logic;
            trigger2      : out std_logic;
            trigger1      : out std_logic;
            pronto_medir2 : out std_logic;
            pronto_medir1 : out std_logic;
            sseg1         : out std_logic_vector(6 downto 0);
            sseg2         : out std_logic_vector(6 downto 0);
            sseg3         : out std_logic_vector(6 downto 0);
            sseg4         : out std_logic_vector(6 downto 0);
            saida_serial  : out std_logic;
            pronto_tx     : out std_logic;
            fim_timer1    : out std_logic;
            fim_timer2    : out std_logic;
            mao_presente  : out std_logic
        );
    end component;

    component hex7seg is
        port (
            hexa : in  std_logic_vector(3 downto 0);
            sseg : out std_logic_vector(6 downto 0)
        );
    end component;

    signal s_pronto_medir1, s_pronto_medir2, s_mao_presente, s_fim_timer1, s_fim_timer2, s_pronto_tx,
           s_zera, s_medir1, s_medir2, s_zera_timer1, s_zera_timer2, s_conta_timer1, s_conta_timer2,
           s_gira_servo, s_partida_tx, s_zera_hc : std_logic;
    
    signal s_db_estado : std_logic_vector(3 downto 0);
	 signal s_sel : std_logic_vector(1 downto 0);
    
begin

    UC: soapga_uc
        port map(
            clock           => clock,
            reset           => reset,
            ligar           => ligar,
            pronto_medir1   => s_pronto_medir1, 
            pronto_medir2   => s_pronto_medir2,
            mao_presente    => s_mao_presente,
            fim_timer1      => s_fim_timer1,
            fim_timer2      => s_fim_timer2,
            pronto_tx       => s_pronto_tx,
            zera            => s_zera,
            medir1          => s_medir1,
            medir2          => s_medir2,
            zera_timer1     => s_zera_timer1,
            zera_timer2     => s_zera_timer2,
            zera_hc         => s_zera_hc,
            conta_timer1    => s_conta_timer1,
            conta_timer2    => s_conta_timer2,
            gira_servo      => s_gira_servo,
            partida_tx      => s_partida_tx,
            sel             => s_sel,
            db_estado       => s_db_estado
        );

    FD: soapga_fd
        port map(
            clock         => clock,
            reset         => s_zera,
            gira_servo    => s_gira_servo,
            medir2        => s_medir2,
            medir1        => s_medir1,
            echo2         => echo2,
            echo1         => echo1,
            sel           => s_sel,
            partida_tx    => s_partida_tx,
            zera_timer1   => s_zera_timer1,
            zera_timer2   => s_zera_timer2,
            zera_hc       => s_zera_hc,
            conta_timer1  => s_conta_timer1,
            conta_timer2  => s_conta_timer2,
            pwm           => pwm,
            trigger2      => trigger2,
            trigger1      => trigger1,
            pronto_medir2 => s_pronto_medir2,
            pronto_medir1 => s_pronto_medir1,
            sseg1         => sseg1,
            sseg2         => sseg2,
            sseg3         => sseg3,
            sseg4         => sseg4,
            saida_serial  => saida_serial,
            pronto_tx     => s_pronto_tx,
            fim_timer1    => s_fim_timer1,
            fim_timer2    => s_fim_timer2,
            mao_presente  => s_mao_presente
        );

    UCSTATE: hex7seg
        port map(
            hexa => s_db_estado,
            sseg => db_estado
        );
        

end architecture;

